��  CCircuit��  CSerializeHack           ��  CPart  (  (      ��� 	 CLogicOut�� 	 CTerminal  �x��      n          �            x���          ��    �
�  �x��               @            ����         ��    �
�  x	�      	         @             ��         ��    �
�  �x��               @            ����         ��    �
�  �x��                �            ����          ��    ��  CLogicIn�� 	 CLatchKey  �a �o          
�  �l ��                             �d �l         ����     ��  �q �         
�  �| ��               @            �t �|        ����     ��  CAND
�  �p�q               �          
�  �`�a              @          
�  �h�i               �            �\�t          ��    ��  CXOR
�  ��                �          
�   ��               @          
�  �	�     	         @            ���    #      ��    �
�  dxyy              @          
�  dhyi                          
�  8pMq               �            Ldd|    '      ��    !�
�  ����                           
�  ����               @          
�  ��)              @            ���    +      ��    �
�  t� ��               @          
�  t� ��               @          
�  H� ]�      k         @            \� t�     /      ��    �
�  �� ��                           
�  �� ��               @          
�  �� ��                �            �� ��     3      ��    �
�  D� Y�      f                     
�  D� Y�      f                     
�  � -�      h          �            ,� D�     7      ��    !�
�  � �      g                     
�  � �      f                     
�  �,�A     i          �            ��,    ;      ��    !�
�  ����               @          
�  ����      i          �          
�  ����              @            ����    ?      ��    ��  COR
�  � �!     j          �          
�  ��     h          �          
�  ��     n          �            ��$    D      ��    �
�  Lpaq              @          
�  L`aa     i          �          
�   h5i     j          �            4\Lt    H      ��    ��  �Y �g       K   
�  �d �y      g                       �\ �d     M    ����     ��  xi �w       N   
�  �t ��      f                       �l �t     P    ����     B�
�   !!               �          
�  !     k         @          
�  ��              @            �$    R      ��    !�
�  ����                �          
�  ����                �          
�  ����               �            ����    V      ��    �
�  tp�q               �          
�  t`�a               �          
�  Hh]i               �            \\tt    Z      ��    !�
�  �� �               @          
�  �� �               @          
�  �$�9               �            ��$    ^      ��    ��  �Y �g      a   
�  �d �y               @            �\ �d     c   ����     ��  �i �w      d   
�  �t ��               @            �l �t     f   ����     ��  �i �w       g   
�  �t ��                             �l �t     i    ����     ��  �Y  g      j   
�  d 	y               @            \ d     l   ����     B�
�  4 I!               �          
�  4I               �          
�                 �            4$    n      ��    !�
�  � 	               @          
�  �� �                           
�   $9              @            �$    r      ��      (  (      ���  CWire  �(�y       v�  �	y      	 v�  ���y       v�  ���y       v�  ��y      n v�  ��     n v�  �@�a      i v�  �       h v�  X� ��      f v�  �p	q      v�  �p�q      v�  Hh�i      v�   hIi      v�   � !      k v�   � I�      k v�  p9q      v�  H Ii       v�  �`a      v�   8a       v��� 
 CCrossOver  �lt         `�       v�  p�       v���  �lt        �pq      v���  �d�l        xh�i      v�  �� �i       v���  �d�l        �� �y       v�  �h��       v�  xx�y      v�  �x��       v�  � �i      j v�  �     h v�  �� ��       f v�  �� �      f v�  X� ��      f v�  �� ��       f v�  �� ��       v���  �� ��         �� ��        v�  �� ��        v���  �� ��         �� ��       v�  �x ��        v�  �� ��        v�  H� I       v�  H� ��       v���  �� ��         �� 	�       v�  x 	�        v���  �� ��         �� ��        v�  � 	�        v�  �� ��       v�  �� ��        v�  �p��       v���  �l�t        `p�q      v�  ``�a     i v���  �l�t        �`��      i v�  ��q       v�  �x �      g v�  �h!i     j v�    !i       v�  �p��       v���  �l�t        �`��       v�  	q       v�  �8�a       v�  �`�a      v���  �l�t        �p�q        (  (      �  (  (        (  (       {   z   x   w   y    �   �   �   �   �   # � # $ � $ % % x ' ' � ( ( � ) � ) + � + , � , - - w / / � 0 0 � 1 � 1 3 3 � 4 4 � 5 � 5 7 7  8 8 � 9 ~ 9 ; � ; < � < = = } ? � ? @ � @ A A z D D � E E � F | F H H � I I � J � J M M � P P � R R � S S � T � T V � V W � W X X y Z Z � [ [ � \ � \ ^ � ^ _ � _ ` ` � c c � f f � i i � l l � n n � o o � p � p r � r s � s t t � -  %  X  A  |  { F = � 9 � 7 � � � � � �   � \ � S � 1 � ) n �  � t � � � � $ � # � �  � � � ( �  � � �  � � + ' � � , D � E ~ �  � < 8 � P � / � � � f � � _ � � 0 � c � � ^ � o � 5 � � 4 � l � � � i � � r 3 � � s � ? � � H � I � � � } @ T � M ; � J R � � V � � � W p � ` � [ � � � Z �  o           �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 